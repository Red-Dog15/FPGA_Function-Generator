
--	 Main Function_Generator File --

--entitiy