-- Button incrementer